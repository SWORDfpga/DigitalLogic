`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:19:38 07/17/2012 
// Design Name: 
// Module Name:    clk_div 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module  clkdiv(input clk,
					output reg[31:0]clkdiv
					);
					
// Clock divider-ʱ�ӷ�Ƶ��

	always @ (posedge clk ) begin 
		clkdiv <= clkdiv + 1'b1; 
	end
	
endmodule
